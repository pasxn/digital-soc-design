library verilog;
use verilog.vl_types.all;
entity mux_2to1_vlg_check_tst is
    port(
        m               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux_2to1_vlg_check_tst;
