library verilog;
use verilog.vl_types.all;
entity andgate_tb is
end andgate_tb;
