library verilog;
use verilog.vl_types.all;
entity mux_5to1_vlg_vec_tst is
end mux_5to1_vlg_vec_tst;
