library verilog;
use verilog.vl_types.all;
entity part_5_vlg_vec_tst is
end part_5_vlg_vec_tst;
