library verilog;
use verilog.vl_types.all;
entity andgate_vlg_check_tst is
    port(
        c               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end andgate_vlg_check_tst;
