library verilog;
use verilog.vl_types.all;
entity seven_segment_decoder_vlg_vec_tst is
end seven_segment_decoder_vlg_vec_tst;
