library verilog;
use verilog.vl_types.all;
entity andgate_vlg_vec_tst is
end andgate_vlg_vec_tst;
